----------------------------------------------------------------------
---------------------//Memory 16 X 16 X 162BitData//--------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.std_logic_arith.all;

entity Memory is
  port(
      Clock: in std_logic;
      Address: in std_logic_vector(7 downto 0);--Address
      Data:in std_logic_vector(162 downto 0);--Always from Accumulator      
      MemEnable:in std_logic;
      RW:in std_logic;
      Output:out std_logic_vector(170 downto 0)
      );
end Memory;
 
architecture Operation of Memory is

begin
  process(Clock)
    type ram is array (0 to 255)of std_logic_vector(170 downto 0);
    variable r:ram;

    begin

   			--write the program here
      --MVI Data
      r(0):="000001000111111000011101011101010010110001010000110101000101101110101111110101000000000000100010001011010001101010010011001010000000000011111101000001101000011111000110110";      
      --MOV Px,A
      r(1):="000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data
      r(2):="000001000000000000000000000001111000110110001110001101000000000100100101111101000101000000010000001000000000000000000000000000000000000111100000000000000000000100111010001";      
      --MOV Py,A
      r(3):="000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";            
      --MVI Data
      r(4):="000001000111111000011101011101000010110001010000110101000101101010101111110101000001001100100010001011010001101010010011001010001100011011111101000001101000011111000110110";      
      --MOV Qx,A
      r(5):="000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data
      r(6):="000001000001101010100011111101111000110110001110001101000000000100100101111101000101100110111010101010001011011000100011100010111000000110001111001011100110010010011110001";      
      --MOV Qy,A
      r(7):="000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data
      r(8):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      --MOV Qz,A
      r(9):="000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 3
	--MUL A,Px
      r(10):="010100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(11):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 4
	--SQR Qz
      r(12):="010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(13):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 5
	--MOV A,T1
      r(14):="000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";     
      --ADD A,Qx
      r(15):="001011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";       
      --MOV X3,A
      r(16):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 6
	--MUL A,Qz
      r(17):="010101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A            
      r(18):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 7
	--MOV A,Py
      r(19):="000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MUL A,T2
      r(20):="010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      --MOV T3,A
      r(21):="000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 8
	--ADD A,Qy
      r(22):="001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(23):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 9
	--MOV A,X3
      r(24):="000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --JZ Address
      r(25):="011010101000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 10
	--SQR A,T1
      r(26):="001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Z3,A
      r(27):="000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 11
	--MOV A,T1
      r(28):="000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MUL A,Y3
      r(29):="010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T3,A      
      r(30):="000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 12
	--MOV A,T1
      r(31):="000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,T2
      r(32):="000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(33):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 13
	--SQR A,X3
      r(34):="001101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(35):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 14
	--MUL A,T1
      r(36):="010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV X3,A
      r(37):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 15
	--SQR A,Y3
      r(38):="001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010001110000";      
      --MOV T2,A
      r(39):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 16
	--ADD A,X3
      r(40):="001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000110000001000000010000010";      
      --MOV X3,A
      r(41):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 17
	--ADD A,T3
      r(42):="000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010001110000";      
      --MOV X3,A
      r(43):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 18
	--MOV A,Px
      r(44):="000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000110000001000000010000010";      
      --MUL A,Z3
      r(45):="010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(46):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000101110010001000000101001000000100000010000000001000";      
      
	--Step 19
	--ADD A,X3
      r(47):="001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(48):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 20
	--SQR A,Z3
      r(49):="001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(50):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 21
	--MOV A,Z3
      r(51):="000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,T3
      r(52):="000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";     
      --MOV T3,A
      r(53):="000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";       
      
	--Step 22
	--MUL A,T2
      r(54):="010010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(55):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 23
	--MOV A,Px          
      r(56):="000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,Py
      r(57):="001010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(58):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      
	--Step 24
	--MUL A,T1
      r(59):="010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T3,A
      r(60):="000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 25
	--ADD A,Y3
      r(61):="001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(62):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Halt
      r(63):="011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(64):="011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      
      --Step 9.1
      --MOV A,Y3
      r(70):="000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";            
      --JZ Address
      r(71):="011010100101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      
	--Step 9.2 if Y3=0
	--MVI Data
      r(72):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      --MOV X3,A
      r(73):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data
      r(74):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(75):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";            
      --MVI Data
      r(76):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Z3,A
      r(77):="000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --Halt
      r(78):="011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      
	--Step 9.1 if Y3=0
      --Point Doubling
      --MOV A,Px
      r(90):="000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Qx,A
      r(91):="000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV A,Py
      r(92):="000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Qy,A
      r(93):="000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data
      r(94):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      --MOV Qz,A
      r(95):="000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --SQR Qz
      r(96):="010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(97):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --SQR Qx
      r(98):="010000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(99):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MUL A,T1
      r(100):="010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";     
      --MOV Z3,A
      r(101):="000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";       
      --SQR T2
      r(102):="001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV X3,A
      r(103):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --SQR T1            
      r(104):="001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(105):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MVI Data(b)
      r(106):="000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";      
      --MUL A,T1
      r(107):="010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T2,A
      r(108):="000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,X3
      r(109):="001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV X3,A
      r(110):="000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --SQR Qy
      r(111):="010001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --Mov T1,A
      r(112):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,Z3
      r(113):="001001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(114):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --ADD A,T2
      r(115):="000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A      
      r(116):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MUL A,X3
      r(117):="010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(118):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV A,T2
      r(119):="000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --NOP
      r(120):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      --MUL A,Z3
      r(121):="010100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV T1,A
      r(122):="000101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --Add A,Y3
      r(123):="001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --MOV Y3,A
      r(124):="000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";      
      --Halt
      r(125):="011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";



      if(MemEnable='1' and Clock='1' and RW='0')then    --Write Operation
        r(conv_integer(Address)):= "00000000" & Data;
      elsif(MemEnable='1' and Clock='1' and RW='1')then --Read Operation 
        Output<=r(conv_integer(Address));
      end if;
    end process;
end Operation;

----------------------------------------------------------------------