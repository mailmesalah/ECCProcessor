----------------------------------------------------------------------
---------------------//Memory 16 X 16 X 162BitData//--------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.std_logic_arith.all;

entity Memory is
  port(
      Clock: in std_logic;
      Address: in std_logic_vector(7 downto 0);--Address
      Data:in std_logic_vector(162 downto 0);--Always from Accumulator      
      MemEnable:in std_logic;
      RW:in std_logic;
      Output:out std_logic_vector(170 downto 0)
      );
end Memory;
 
architecture Operation of Memory is

begin
  process(Clock)
    type ram is array (0 to 255)of std_logic_vector(170 downto 0);
    variable r:ram;

    begin
      --write the program here
      r(0):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(1):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(2):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(3):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(4):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
      r(5):="000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

      if(MemEnable='1' and Clock='1' and RW='0')then    --Write Operation
        r(conv_integer(Address)):= "00000000" & Data;
      elsif(MemEnable='1' and Clock='1' and RW='1')then --Read Operation 
        Output<=r(conv_integer(Address));
      end if;
    end process;
end Operation;

----------------------------------------------------------------------