----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:44:14 07/15/2013 
-- Design Name: 
-- Module Name:    full_163bitmul - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Mul is
    Port( 
        a : in  STD_LOGIC_VECTOR (162 downto 0);
        b : in  STD_LOGIC;
        clk : in  STD_LOGIC;
        reset : in  STD_LOGIC;
        c : out  STD_LOGIC_VECTOR (162 downto 0));
end Mul;

architecture Behavioral of Mul is
   signal sig_0  : std_logic;
   signal sig_1  : std_logic;
   signal sig_2  : std_logic;
   signal sig_3  : std_logic;
   signal sig_4  : std_logic;
   signal sig_5  : std_logic;
   signal sig_6  : std_logic;
   signal sig_7  : std_logic;
   signal sig_8  : std_logic;
   signal sig_9  : std_logic;
   signal sig_10 : std_logic;
   signal sig_11 : std_logic;
   signal sig_12 : std_logic;
   signal sig_13 : std_logic;
   signal sig_14 : std_logic;
   signal sig_15 : std_logic;
   signal sig_16 : std_logic;
   signal sig_17 : std_logic;
   signal sig_18 : std_logic;
   signal sig_19 : std_logic;
   signal sig_20 : std_logic;
   signal sig_21 : std_logic;
   signal sig_22 : std_logic;
   signal sig_23 : std_logic;
   signal sig_24 : std_logic;
   signal sig_25 : std_logic;
   signal sig_26 : std_logic;
   signal sig_27 : std_logic;
   signal sig_28 : std_logic;
   signal sig_29 : std_logic;
   signal sig_30 : std_logic;
   signal sig_31 : std_logic;
   signal sig_32 : std_logic;
   signal sig_33 : std_logic;
   signal sig_34 : std_logic;
   signal sig_35 : std_logic;
   signal sig_36 : std_logic;
   signal sig_37 : std_logic;
   signal sig_38 : std_logic;
   signal sig_39 : std_logic;
   signal sig_40 : std_logic;
   signal sig_41 : std_logic;
   signal sig_42 : std_logic;
   signal sig_43 : std_logic;
   signal sig_44 : std_logic;
   signal sig_45 : std_logic;
   signal sig_46 : std_logic;
   signal sig_47 : std_logic;
   signal sig_48 : std_logic;
   signal sig_49 : std_logic;
   signal sig_50 : std_logic;
   signal sig_51 : std_logic;
   signal sig_52 : std_logic;
   signal sig_53 : std_logic;
   signal sig_54 : std_logic;
   signal sig_55 : std_logic;
   signal sig_56 : std_logic;
   signal sig_57 : std_logic;
   signal sig_58 : std_logic;
   signal sig_59 : std_logic;
   signal sig_60 : std_logic;
   signal sig_61 : std_logic;
   signal sig_62 : std_logic;
   signal sig_63 : std_logic;
   signal sig_64 : std_logic;
   signal sig_65 : std_logic;
   signal sig_66 : std_logic;
   signal sig_67 : std_logic;
   signal sig_68 : std_logic;
   signal sig_69 : std_logic;
   signal sig_70 : std_logic;
   signal sig_71 : std_logic;
   signal sig_72 : std_logic;
   signal sig_73 : std_logic;
   signal sig_74 : std_logic;
   signal sig_75 : std_logic;
   signal sig_76 : std_logic;
   signal sig_77 : std_logic;
   signal sig_78 : std_logic;
   signal sig_79 : std_logic;
   signal sig_80 : std_logic;
   signal sig_81 : std_logic;
   signal sig_82 : std_logic;
   signal sig_83 : std_logic;
   signal sig_84 : std_logic;
   signal sig_85 : std_logic;
   signal sig_86 : std_logic;
   signal sig_87 : std_logic;
   signal sig_88 : std_logic;
   signal sig_89 : std_logic;
   signal sig_90 : std_logic;
   signal sig_91 : std_logic;
   signal sig_92 : std_logic;
   signal sig_93 : std_logic;
   signal sig_94 : std_logic;
   signal sig_95 : std_logic;
   signal sig_96 : std_logic;
   signal sig_97 : std_logic;
   signal sig_98 : std_logic;
   signal sig_99 : std_logic;
   signal sig_100: std_logic;
   signal sig_101: std_logic;
   signal sig_102: std_logic;
   signal sig_103: std_logic;
   signal sig_104: std_logic;
   signal sig_105: std_logic;
   signal sig_106: std_logic;
   signal sig_107: std_logic;
   signal sig_108: std_logic;
   signal sig_109: std_logic;
   signal sig_110: std_logic;
   signal sig_111: std_logic;
   signal sig_112: std_logic;
   signal sig_113: std_logic;
   signal sig_114: std_logic;
   signal sig_115: std_logic;
   signal sig_116: std_logic;
   signal sig_117: std_logic;
   signal sig_118: std_logic;
   signal sig_119: std_logic;
   signal sig_120: std_logic;
   signal sig_121: std_logic;
   signal sig_122: std_logic;
   signal sig_123: std_logic;
   signal sig_124: std_logic;
   signal sig_125: std_logic;
   signal sig_126: std_logic;
   signal sig_127: std_logic;
   signal sig_128: std_logic;
   signal sig_129: std_logic;
   signal sig_130: std_logic;
   signal sig_131: std_logic;
   signal sig_132: std_logic;
   signal sig_133: std_logic;
   signal sig_134: std_logic;
   signal sig_135: std_logic;
   signal sig_136: std_logic;
   signal sig_137: std_logic;
   signal sig_138: std_logic;
   signal sig_139: std_logic;
   signal sig_140: std_logic;
   signal sig_141: std_logic;
   signal sig_142: std_logic;
   signal sig_143: std_logic;
   signal sig_144: std_logic;
   signal sig_145: std_logic;
   signal sig_146: std_logic;
   signal sig_147: std_logic;
   signal sig_148: std_logic;
   signal sig_149: std_logic;
   signal sig_150: std_logic;
   signal sig_151: std_logic;
   signal sig_152: std_logic;
   signal sig_153: std_logic;
   signal sig_154: std_logic;
   signal sig_155: std_logic;
   signal sig_156: std_logic;
   signal sig_157: std_logic;
   signal sig_158: std_logic;
   signal sig_159: std_logic;
   signal sig_160: std_logic;
   signal sig_161: std_logic;
   signal sig_162: std_logic;
   signal xor_0     : std_logic;
   signal xor_1     : std_logic;
   signal xor_2     : std_logic;
   signal xor_3     : std_logic;
   signal xor_4     : std_logic;
   signal xor_5     : std_logic;
   signal xor_6     : std_logic;
   signal xor_7     : std_logic;
   signal xor_8     : std_logic;
   signal xor_9     : std_logic;
   signal xor_10    : std_logic;
   signal xor_11    : std_logic;
   signal xor_12    : std_logic;
   signal xor_13    : std_logic;
   signal xor_14    : std_logic;
   signal xor_15    : std_logic;
   signal xor_16    : std_logic;
   signal xor_17    : std_logic;
   signal xor_18    : std_logic;
   signal xor_19    : std_logic;
   signal xor_20    : std_logic;
   signal xor_21    : std_logic;
   signal xor_22    : std_logic;
   signal xor_23    : std_logic;
   signal xor_24    : std_logic;
   signal xor_25    : std_logic;
   signal xor_26    : std_logic;
   signal xor_27    : std_logic;
   signal xor_28    : std_logic;
   signal xor_29    : std_logic;
   signal xor_30    : std_logic;
   signal xor_31    : std_logic;
   signal xor_32    : std_logic;
   signal xor_33    : std_logic;
   signal xor_34    : std_logic;
   signal xor_35    : std_logic;
   signal xor_36    : std_logic;
   signal xor_37    : std_logic;
   signal xor_38    : std_logic;
   signal xor_39    : std_logic;
   signal xor_40    : std_logic;
   signal xor_41    : std_logic;
   signal xor_42    : std_logic;
   signal xor_43    : std_logic;
   signal xor_44    : std_logic;
   signal xor_45    : std_logic;
   signal xor_46    : std_logic;
   signal xor_47    : std_logic;
   signal xor_48    : std_logic;
   signal xor_49    : std_logic;
   signal xor_50    : std_logic;
   signal xor_51    : std_logic;
   signal xor_52    : std_logic;
   signal xor_53    : std_logic;
   signal xor_54    : std_logic;
   signal xor_55    : std_logic;
   signal xor_56    : std_logic;
   signal xor_57    : std_logic;
   signal xor_58    : std_logic;
   signal xor_59    : std_logic;
   signal xor_60    : std_logic;
   signal xor_61    : std_logic;
   signal xor_62    : std_logic;
   signal xor_63    : std_logic;
   signal xor_64    : std_logic;
   signal xor_65    : std_logic;
   signal xor_66    : std_logic;
   signal xor_67    : std_logic;
   signal xor_68    : std_logic;
   signal xor_69    : std_logic;
   signal xor_70    : std_logic;
   signal xor_71    : std_logic;
   signal xor_72    : std_logic;
   signal xor_73    : std_logic;
   signal xor_74    : std_logic;
   signal xor_75    : std_logic;
   signal xor_76    : std_logic;
   signal xor_77    : std_logic;
   signal xor_78    : std_logic;
   signal xor_79    : std_logic;
   signal xor_80    : std_logic;
   signal xor_81    : std_logic;
   signal xor_82    : std_logic;
   signal xor_83    : std_logic;
   signal xor_84    : std_logic;
   signal xor_85    : std_logic;
   signal xor_86    : std_logic;
   signal xor_87    : std_logic;
   signal xor_88    : std_logic;
   signal xor_89    : std_logic;
   signal xor_90    : std_logic;
   signal xor_91    : std_logic;
   signal xor_92    : std_logic;
   signal xor_93    : std_logic;
   signal xor_94    : std_logic;
   signal xor_95    : std_logic;
   signal xor_96    : std_logic;
   signal xor_97    : std_logic;
   signal xor_98    : std_logic;
   signal xor_99    : std_logic;
   signal xor_100   : std_logic;
   signal xor_101   : std_logic;
   signal xor_102   : std_logic;
   signal xor_103   : std_logic;
   signal xor_104   : std_logic;
   signal xor_105   : std_logic;
   signal xor_106   : std_logic;
   signal xor_107   : std_logic;
   signal xor_108   : std_logic;
   signal xor_109   : std_logic;
   signal xor_110   : std_logic;
   signal xor_111   : std_logic;
   signal xor_112   : std_logic;
   signal xor_113   : std_logic;
   signal xor_114   : std_logic;
   signal xor_115   : std_logic;
   signal xor_116   : std_logic;
   signal xor_117   : std_logic;
   signal xor_118   : std_logic;
   signal xor_119   : std_logic;
   signal xor_120   : std_logic;
   signal xor_121   : std_logic;
   signal xor_122   : std_logic;
   signal xor_123   : std_logic;
   signal xor_124   : std_logic;
   signal xor_125   : std_logic;
   signal xor_126   : std_logic;
   signal xor_127   : std_logic;
   signal xor_128   : std_logic;
   signal xor_129   : std_logic;
   signal xor_130   : std_logic;
   signal xor_131   : std_logic;
   signal xor_132   : std_logic;
   signal xor_133   : std_logic;
   signal xor_134   : std_logic;
   signal xor_135   : std_logic;
   signal xor_136   : std_logic;
   signal xor_137   : std_logic;
   signal xor_138   : std_logic;
   signal xor_139   : std_logic;
   signal xor_140   : std_logic;
   signal xor_141   : std_logic;
   signal xor_142   : std_logic;
   signal xor_143   : std_logic;
   signal xor_144   : std_logic;
   signal xor_145   : std_logic;
   signal xor_146   : std_logic;
   signal xor_147   : std_logic;
   signal xor_148   : std_logic;
   signal xor_149   : std_logic;
   signal xor_150   : std_logic;
   signal xor_151   : std_logic;
   signal xor_152   : std_logic;
   signal xor_153   : std_logic;
   signal xor_154   : std_logic;
   signal xor_155   : std_logic;
   signal xor_156   : std_logic;
   signal xor_157   : std_logic;
   signal xor_158   : std_logic;
   signal xor_159   : std_logic;
   signal xor_160   : std_logic;
   signal xor_161   : std_logic;
   signal xor_162   : std_logic;
   signal c0_DUMMY  : std_logic;
   signal c1_DUMMY  : std_logic;
   signal c2_DUMMY  : std_logic;
   signal c3_DUMMY  : std_logic;
   signal c4_DUMMY  : std_logic;
   signal c5_DUMMY  : std_logic;
   signal c6_DUMMY  : std_logic;
   signal c7_DUMMY  : std_logic;
   signal c8_DUMMY  : std_logic;
   signal c9_DUMMY  : std_logic;
   signal c10_DUMMY  : std_logic;
   signal c11_DUMMY  : std_logic;
   signal c12_DUMMY  : std_logic;
   signal c13_DUMMY  : std_logic;
   signal c14_DUMMY  : std_logic;
   signal c15_DUMMY  : std_logic;
   signal c16_DUMMY  : std_logic;
   signal c17_DUMMY  : std_logic;
   signal c18_DUMMY  : std_logic;
   signal c19_DUMMY  : std_logic;
   signal c20_DUMMY  : std_logic;
   signal c21_DUMMY  : std_logic;
   signal c22_DUMMY  : std_logic;
   signal c23_DUMMY  : std_logic;
   signal c24_DUMMY  : std_logic;
   signal c25_DUMMY  : std_logic;
   signal c26_DUMMY  : std_logic;
   signal c27_DUMMY  : std_logic;
   signal c28_DUMMY  : std_logic;
   signal c29_DUMMY  : std_logic;
   signal c30_DUMMY  : std_logic;
   signal c31_DUMMY  : std_logic;
   signal c32_DUMMY  : std_logic;
   signal c33_DUMMY  : std_logic;
   signal c34_DUMMY  : std_logic;
   signal c35_DUMMY  : std_logic;
   signal c36_DUMMY  : std_logic;
   signal c37_DUMMY  : std_logic;
   signal c38_DUMMY  : std_logic;
   signal c39_DUMMY  : std_logic;
   signal c40_DUMMY  : std_logic;
   signal c41_DUMMY  : std_logic;
   signal c42_DUMMY  : std_logic;
   signal c43_DUMMY  : std_logic;
   signal c44_DUMMY  : std_logic;
   signal c45_DUMMY  : std_logic;
   signal c46_DUMMY  : std_logic;
   signal c47_DUMMY  : std_logic;
   signal c48_DUMMY  : std_logic;
   signal c49_DUMMY  : std_logic;
   signal c50_DUMMY  : std_logic;
   signal c51_DUMMY  : std_logic;
   signal c52_DUMMY  : std_logic;
   signal c53_DUMMY  : std_logic;
   signal c54_DUMMY  : std_logic;
   signal c55_DUMMY  : std_logic;
   signal c56_DUMMY  : std_logic;
   signal c57_DUMMY  : std_logic;
   signal c58_DUMMY  : std_logic;
   signal c59_DUMMY  : std_logic;
   signal c60_DUMMY  : std_logic;
   signal c61_DUMMY  : std_logic;
   signal c62_DUMMY  : std_logic;
   signal c63_DUMMY  : std_logic;
   signal c64_DUMMY  : std_logic;
   signal c65_DUMMY  : std_logic;
   signal c66_DUMMY  : std_logic;
   signal c67_DUMMY  : std_logic;
   signal c68_DUMMY  : std_logic;
   signal c69_DUMMY  : std_logic;
   signal c70_DUMMY  : std_logic;
   signal c71_DUMMY  : std_logic;
   signal c72_DUMMY  : std_logic;
   signal c73_DUMMY  : std_logic;
   signal c74_DUMMY  : std_logic;
   signal c75_DUMMY  : std_logic;
   signal c76_DUMMY  : std_logic;
   signal c77_DUMMY  : std_logic;
   signal c78_DUMMY  : std_logic;
   signal c79_DUMMY  : std_logic;
   signal c80_DUMMY  : std_logic;
   signal c81_DUMMY  : std_logic;
   signal c82_DUMMY  : std_logic;
   signal c83_DUMMY  : std_logic;
   signal c84_DUMMY  : std_logic;
   signal c85_DUMMY  : std_logic;
   signal c86_DUMMY  : std_logic;
   signal c87_DUMMY  : std_logic;
   signal c88_DUMMY  : std_logic;
   signal c89_DUMMY  : std_logic;
   signal c90_DUMMY  : std_logic;
   signal c91_DUMMY  : std_logic;
   signal c92_DUMMY  : std_logic;
   signal c93_DUMMY  : std_logic;
   signal c94_DUMMY  : std_logic;
   signal c95_DUMMY  : std_logic;
   signal c96_DUMMY  : std_logic;
   signal c97_DUMMY  : std_logic;
   signal c98_DUMMY  : std_logic;
   signal c99_DUMMY  : std_logic;
   signal c100_DUMMY  : std_logic;
   signal c101_DUMMY  : std_logic;
   signal c102_DUMMY  : std_logic;
   signal c103_DUMMY  : std_logic;
   signal c104_DUMMY  : std_logic;
   signal c105_DUMMY  : std_logic;
   signal c106_DUMMY  : std_logic;
   signal c107_DUMMY  : std_logic;
   signal c108_DUMMY  : std_logic;
   signal c109_DUMMY  : std_logic;
   signal c110_DUMMY  : std_logic;
   signal c111_DUMMY  : std_logic;
   signal c112_DUMMY  : std_logic;
   signal c113_DUMMY  : std_logic;
   signal c114_DUMMY  : std_logic;
   signal c115_DUMMY  : std_logic;
   signal c116_DUMMY  : std_logic;
   signal c117_DUMMY  : std_logic;
   signal c118_DUMMY  : std_logic;
   signal c119_DUMMY  : std_logic;
   signal c120_DUMMY  : std_logic;
   signal c121_DUMMY  : std_logic;
   signal c122_DUMMY  : std_logic;
   signal c123_DUMMY  : std_logic;
   signal c124_DUMMY  : std_logic;
   signal c125_DUMMY  : std_logic;
   signal c126_DUMMY  : std_logic;
   signal c127_DUMMY  : std_logic;
   signal c128_DUMMY  : std_logic;
   signal c129_DUMMY  : std_logic;
   signal c130_DUMMY  : std_logic;
   signal c131_DUMMY  : std_logic;
   signal c132_DUMMY  : std_logic;
   signal c133_DUMMY  : std_logic;
   signal c134_DUMMY  : std_logic;
   signal c135_DUMMY  : std_logic;
   signal c136_DUMMY  : std_logic;
   signal c137_DUMMY  : std_logic;
   signal c138_DUMMY  : std_logic;
   signal c139_DUMMY  : std_logic;
   signal c140_DUMMY  : std_logic;
   signal c141_DUMMY  : std_logic;
   signal c142_DUMMY  : std_logic;
   signal c143_DUMMY  : std_logic;
   signal c144_DUMMY  : std_logic;
   signal c145_DUMMY  : std_logic;
   signal c146_DUMMY  : std_logic;
   signal c147_DUMMY  : std_logic;
   signal c148_DUMMY  : std_logic;
   signal c149_DUMMY  : std_logic;
   signal c150_DUMMY  : std_logic;
   signal c151_DUMMY  : std_logic;
   signal c152_DUMMY  : std_logic;
   signal c153_DUMMY  : std_logic;
   signal c154_DUMMY  : std_logic;
   signal c155_DUMMY  : std_logic;
   signal c156_DUMMY  : std_logic;
   signal c157_DUMMY  : std_logic;
   signal c158_DUMMY  : std_logic;
   signal c159_DUMMY  : std_logic;
   signal c160_DUMMY  : std_logic;
   signal c161_DUMMY  : std_logic;
   signal c162_DUMMY  : std_logic;
   signal xor_c2c162  : std_logic;
   signal xor_c5c162  : std_logic;
   signal xor_c6c162  : std_logic;
component and_2
port ( I0 : in    std_logic; 
       I1 : in    std_logic; 
       o  : out   std_logic);
   end component;
component xor_2b
      port ( I0 : in    std_logic; 
             I1 : in    std_logic; 
             o  : out   std_logic);
   end component;
component reg_dff
      port (  D : in    std_logic; 
             clk : in    std_logic;
             reset : in std_logic;			 
             Q : out   std_logic);
	end component;	

begin
sigI_0 : and_2
      port map (I0=>a(0),
                I1=>b,
                O=>sig_0);
sigI_1 : and_2
      port map (I0=>a(1),
                I1=>b,
                O=>sig_1);
sigI_2 : and_2
      port map (I0=>a(2),
                I1=>b,
                O=>sig_2);
sigI_3 : and_2
      port map (I0=>a(3),
                I1=>b,
                O=>sig_3);
sigI_4 : and_2
      port map (I0=>a(4),
                I1=>b,
                O=>sig_4);
sigI_5 : and_2
      port map (I0=>a(5),
                I1=>b,
                O=>sig_5);
sigI_6 : and_2
      port map (I0=>a(6),
                I1=>b,
                O=>sig_6);
sigI_7 : and_2
      port map (I0=>a(7),
                I1=>b,
                O=>sig_7);
sigI_8 : and_2
      port map (I0=>a(8),
                I1=>b,
                O=>sig_8);
sigI_9 : and_2
      port map (I0=>a(9),
                I1=>b,
                O=>sig_9);
sigI_10 : and_2
      port map (I0=>a(10),
                I1=>b,
                O=>sig_10);
sigI_11 : and_2
      port map (I0=>a(11),
                I1=>b,
                O=>sig_11);
sigI_12 : and_2
      port map (I0=>a(12),
                I1=>b,
                O=>sig_12);
sigI_13 : and_2
      port map (I0=>a(13),
                I1=>b,
                O=>sig_13);
sigI_14 : and_2
      port map (I0=>a(14),
                I1=>b,
                O=>sig_14);
sigI_15 : and_2
      port map (I0=>a(15),
                I1=>b,
                O=>sig_15);
sigI_16 : and_2
      port map (I0=>a(16),
                I1=>b,
                O=>sig_16);
sigI_17 : and_2
      port map (I0=>a(17),
                I1=>b,
                O=>sig_17);
sigI_18 : and_2
      port map (I0=>a(18),
                I1=>b,
                O=>sig_18);
sigI_19 : and_2
      port map (I0=>a(19),
                I1=>b,
                O=>sig_19);
sigI_20 : and_2
      port map (I0=>a(20),
                I1=>b,
                O=>sig_20);
sigI_21 : and_2
      port map (I0=>a(21),
                I1=>b,
                O=>sig_21);
sigI_22 : and_2
      port map (I0=>a(22),
                I1=>b,
                O=>sig_22);
sigI_23 : and_2
      port map (I0=>a(23),
                I1=>b,
                O=>sig_23);
sigI_24 : and_2
      port map (I0=>a(24),
                I1=>b,
                O=>sig_24);
sigI_25 : and_2
      port map (I0=>a(25),
                I1=>b,
                O=>sig_25);
sigI_26 : and_2
      port map (I0=>a(26),
                I1=>b,
                O=>sig_26);
sigI_27 : and_2
      port map (I0=>a(27),
                I1=>b,
                O=>sig_27);
sigI_28 : and_2
      port map (I0=>a(28),
                I1=>b,
                O=>sig_28);
sigI_29 : and_2
      port map (I0=>a(29),
                I1=>b,
                O=>sig_29);
sigI_30 : and_2
      port map (I0=>a(30),
                I1=>b,
                O=>sig_30);
sigI_31 : and_2
      port map (I0=>a(31),
                I1=>b,
                O=>sig_31);
sigI_32 : and_2
      port map (I0=>a(32),
                I1=>b,
                O=>sig_32);
sigI_33 : and_2
      port map (I0=>a(33),
                I1=>b,
                O=>sig_33);
sigI_34 : and_2
      port map (I0=>a(34),
                I1=>b,
                O=>sig_34);
sigI_35 : and_2
      port map (I0=>a(35),
                I1=>b,
                O=>sig_35);
sigI_36 : and_2
      port map (I0=>a(36),
                I1=>b,
                O=>sig_36);
sigI_37 : and_2
      port map (I0=>a(37),
                I1=>b,
                O=>sig_37);
sigI_38 : and_2
      port map (I0=>a(38),
                I1=>b,
                O=>sig_38);
sigI_39 : and_2
      port map (I0=>a(39),
                I1=>b,
                O=>sig_39);
sigI_40 : and_2
      port map (I0=>a(40),
                I1=>b,
                O=>sig_40);
sigI_41 : and_2
      port map (I0=>a(41),
                I1=>b,
                O=>sig_41);
sigI_42 : and_2
      port map (I0=>a(42),
                I1=>b,
                O=>sig_42);
sigI_43 : and_2
      port map (I0=>a(43),
                I1=>b,
                O=>sig_43);
sigI_44 : and_2
      port map (I0=>a(44),
                I1=>b,
                O=>sig_44);
sigI_45 : and_2
      port map (I0=>a(45),
                I1=>b,
                O=>sig_45);
sigI_46 : and_2
      port map (I0=>a(46),
                I1=>b,
                O=>sig_46);
sigI_47 : and_2
      port map (I0=>a(47),
                I1=>b,
                O=>sig_47);
sigI_48 : and_2
      port map (I0=>a(48),
                I1=>b,
                O=>sig_48);
sigI_49 : and_2
      port map (I0=>a(49),
                I1=>b,
                O=>sig_49);
sigI_50 : and_2
      port map (I0=>a(50),
                I1=>b,
                O=>sig_50);
sigI_51 : and_2
      port map (I0=>a(51),
                I1=>b,
                O=>sig_51);
sigI_52 : and_2
      port map (I0=>a(52),
                I1=>b,
                O=>sig_52);
sigI_53 : and_2
      port map (I0=>a(53),
                I1=>b,
                O=>sig_53);
sigI_54 : and_2
      port map (I0=>a(54),
                I1=>b,
                O=>sig_54);
sigI_55 : and_2
      port map (I0=>a(55),
                I1=>b,
                O=>sig_55);
sigI_56 : and_2
      port map (I0=>a(56),
                I1=>b,
                O=>sig_56);
sigI_57 : and_2
      port map (I0=>a(57),
                I1=>b,
                O=>sig_57);
sigI_58 : and_2
      port map (I0=>a(58),
                I1=>b,
                O=>sig_58);
sigI_59 : and_2
      port map (I0=>a(59),
                I1=>b,
                O=>sig_59);
sigI_60 : and_2
      port map (I0=>a(60),
                I1=>b,
                O=>sig_60);
sigI_61 : and_2
      port map (I0=>a(61),
                I1=>b,
                O=>sig_61);
sigI_62 : and_2
      port map (I0=>a(62),
                I1=>b,
                O=>sig_62);
sigI_63 : and_2
      port map (I0=>a(63),
                I1=>b,
                O=>sig_63);
sigI_64 : and_2
      port map (I0=>a(64),
                I1=>b,
                O=>sig_64);
sigI_65 : and_2
      port map (I0=>a(65),
                I1=>b,
                O=>sig_65);
sigI_66 : and_2
      port map (I0=>a(66),
                I1=>b,
                O=>sig_66);
sigI_67 : and_2
      port map (I0=>a(67),
                I1=>b,
                O=>sig_67);
sigI_68 : and_2
      port map (I0=>a(68),
                I1=>b,
                O=>sig_68);
sigI_69 : and_2
      port map (I0=>a(69),
                I1=>b,
                O=>sig_69);
sigI_70 : and_2
      port map (I0=>a(70),
                I1=>b,
                O=>sig_70);
sigI_71 : and_2
      port map (I0=>a(71),
                I1=>b,
                O=>sig_71);
sigI_72 : and_2
      port map (I0=>a(72),
                I1=>b,
                O=>sig_72);
sigI_73 : and_2
      port map (I0=>a(73),
                I1=>b,
                O=>sig_73);
sigI_74 : and_2
      port map (I0=>a(74),
                I1=>b,
                O=>sig_74);
sigI_75 : and_2
      port map (I0=>a(75),
                I1=>b,
                O=>sig_75);
sigI_76 : and_2
      port map (I0=>a(76),
                I1=>b,
                O=>sig_76);
sigI_77 : and_2
      port map (I0=>a(77),
                I1=>b,
                O=>sig_77);
sigI_78 : and_2
      port map (I0=>a(78),
                I1=>b,
                O=>sig_78);
sigI_79 : and_2
      port map (I0=>a(79),
                I1=>b,
                O=>sig_79);
sigI_80 : and_2
      port map (I0=>a(80),
                I1=>b,
                O=>sig_80);
sigI_81 : and_2
      port map (I0=>a(81),
                I1=>b,
                O=>sig_81);
sigI_82 : and_2
      port map (I0=>a(82),
                I1=>b,
                O=>sig_82);
sigI_83 : and_2
      port map (I0=>a(83),
                I1=>b,
                O=>sig_83);
sigI_84 : and_2
      port map (I0=>a(84),
                I1=>b,
                O=>sig_84);
sigI_85 : and_2
      port map (I0=>a(85),
                I1=>b,
                O=>sig_85);
sigI_86 : and_2
      port map (I0=>a(86),
                I1=>b,
                O=>sig_86);
sigI_87 : and_2
      port map (I0=>a(87),
                I1=>b,
                O=>sig_87);
sigI_88 : and_2
      port map (I0=>a(88),
                I1=>b,
                O=>sig_88);
sigI_89 : and_2
      port map (I0=>a(89),
                I1=>b,
                O=>sig_89);
sigI_90 : and_2
      port map (I0=>a(90),
                I1=>b,
                O=>sig_90);
sigI_91 : and_2
      port map (I0=>a(91),
                I1=>b,
                O=>sig_91);
sigI_92 : and_2
      port map (I0=>a(92),
                I1=>b,
                O=>sig_92);
sigI_93 : and_2
      port map (I0=>a(93),
                I1=>b,
                O=>sig_93);
sigI_94 : and_2
      port map (I0=>a(94),
                I1=>b,
                O=>sig_94);
sigI_95 : and_2
      port map (I0=>a(95),
                I1=>b,
                O=>sig_95);
sigI_96 : and_2
      port map (I0=>a(96),
                I1=>b,
                O=>sig_96);
sigI_97 : and_2
      port map (I0=>a(97),
                I1=>b,
                O=>sig_97);
sigI_98 : and_2
      port map (I0=>a(98),
                I1=>b,
                O=>sig_98);
sigI_99 : and_2
      port map (I0=>a(99),
                I1=>b,
                O=>sig_99);
sigI_100 : and_2
      port map (I0=>a(100),
                I1=>b,
                O=>sig_100);
sigI_101 : and_2
      port map (I0=>a(101),
                I1=>b,
                O=>sig_101);
sigI_102 : and_2
      port map (I0=>a(102),
                I1=>b,
                O=>sig_102);
sigI_103 : and_2
      port map (I0=>a(103),
                I1=>b,
                O=>sig_103);
sigI_104 : and_2
      port map (I0=>a(104),
                I1=>b,
                O=>sig_104);
sigI_105 : and_2
      port map (I0=>a(105),
                I1=>b,
                O=>sig_105);
sigI_106 : and_2
      port map (I0=>a(106),
                I1=>b,
                O=>sig_106);
sigI_107 : and_2
      port map (I0=>a(107),
                I1=>b,
                O=>sig_107);
sigI_108 : and_2
      port map (I0=>a(108),
                I1=>b,
                O=>sig_108);
sigI_109 : and_2
      port map (I0=>a(109),
                I1=>b,
                O=>sig_109);
sigI_110 : and_2
      port map (I0=>a(110),
                I1=>b,
                O=>sig_110);
sigI_111 : and_2
      port map (I0=>a(111),
                I1=>b,
                O=>sig_111);
sigI_112 : and_2
      port map (I0=>a(112),
                I1=>b,
                O=>sig_112);
sigI_113 : and_2
      port map (I0=>a(113),
                I1=>b,
                O=>sig_113);
sigI_114 : and_2
      port map (I0=>a(114),
                I1=>b,
                O=>sig_114);
sigI_115 : and_2
      port map (I0=>a(115),
                I1=>b,
                O=>sig_115);
sigI_116 : and_2
      port map (I0=>a(116),
                I1=>b,
                O=>sig_116);
sigI_117 : and_2
      port map (I0=>a(117),
                I1=>b,
                O=>sig_117);
sigI_118 : and_2
      port map (I0=>a(118),
                I1=>b,
                O=>sig_118);
sigI_119 : and_2
      port map (I0=>a(119),
                I1=>b,
                O=>sig_119);
sigI_120 : and_2
      port map (I0=>a(120),
                I1=>b,
                O=>sig_120);
sigI_121 : and_2
      port map (I0=>a(121),
                I1=>b,
                O=>sig_121);
sigI_122 : and_2
      port map (I0=>a(122),
                I1=>b,
                O=>sig_122);
sigI_123 : and_2
      port map (I0=>a(123),
                I1=>b,
                O=>sig_123);
sigI_124 : and_2
      port map (I0=>a(124),
                I1=>b,
                O=>sig_124);
sigI_125 : and_2
      port map (I0=>a(125),
                I1=>b,
                O=>sig_125);
sigI_126 : and_2
      port map (I0=>a(126),
                I1=>b,
                O=>sig_126);
sigI_127 : and_2
      port map (I0=>a(127),
                I1=>b,
                O=>sig_127);
sigI_128 : and_2
      port map (I0=>a(128),
                I1=>b,
                O=>sig_128);
sigI_129 : and_2
      port map (I0=>a(129),
                I1=>b,
                O=>sig_129);
sigI_130 : and_2
      port map (I0=>a(130),
                I1=>b,
                O=>sig_130);
sigI_131 : and_2
      port map (I0=>a(131),
                I1=>b,
                O=>sig_131);
sigI_132 : and_2
      port map (I0=>a(132),
                I1=>b,
                O=>sig_132);
sigI_133 : and_2
      port map (I0=>a(133),
                I1=>b,
                O=>sig_133);
sigI_134 : and_2
      port map (I0=>a(134),
                I1=>b,
                O=>sig_134);
sigI_135 : and_2
      port map (I0=>a(135),
                I1=>b,
                O=>sig_135);
sigI_136 : and_2
      port map (I0=>a(136),
                I1=>b,
                O=>sig_136);
sigI_137 : and_2
      port map (I0=>a(137),
                I1=>b,
                O=>sig_137);
sigI_138 : and_2
      port map (I0=>a(138),
                I1=>b,
                O=>sig_138);
sigI_139 : and_2
      port map (I0=>a(139),
                I1=>b,
                O=>sig_139);
sigI_140 : and_2
      port map (I0=>a(140),
                I1=>b,
                O=>sig_140);
sigI_141 : and_2
      port map (I0=>a(141),
                I1=>b,
                O=>sig_141);
sigI_142 : and_2
      port map (I0=>a(142),
                I1=>b,
                O=>sig_142);
sigI_143 : and_2
      port map (I0=>a(143),
                I1=>b,
                O=>sig_143);
sigI_144 : and_2
      port map (I0=>a(144),
                I1=>b,
                O=>sig_144);
sigI_145 : and_2
      port map (I0=>a(145),
                I1=>b,
                O=>sig_145);
sigI_146 : and_2
      port map (I0=>a(146),
                I1=>b,
                O=>sig_146);				
sigI_147 : and_2
      port map (I0=>a(147),
                I1=>b,
                O=>sig_147);
sigI_148 : and_2
      port map (I0=>a(148),
                I1=>b,
                O=>sig_148);
sigI_149 : and_2
      port map (I0=>a(149),
                I1=>b,
                O=>sig_149);
sigI_150 : and_2
      port map (I0=>a(150),
                I1=>b,
                O=>sig_150);
sigI_151 : and_2
      port map (I0=>a(151),
                I1=>b,
                O=>sig_151);
sigI_152 : and_2
      port map (I0=>a(152),
                I1=>b,
                O=>sig_152);
sigI_153 : and_2
      port map (I0=>a(153),
                I1=>b,
                O=>sig_153);
sigI_154 : and_2
      port map (I0=>a(154),
                I1=>b,
                O=>sig_154);
sigI_155 : and_2
      port map (I0=>a(155),
                I1=>b,
                O=>sig_155);
sigI_156 : and_2
      port map (I0=>a(156),
                I1=>b,
                O=>sig_156);
sigI_157 : and_2
      port map (I0=>a(157),
                I1=>b,
                O=>sig_157);
sigI_158 : and_2
      port map (I0=>a(158),
                I1=>b,
                O=>sig_158);
sigI_159 : and_2
      port map (I0=>a(159),
                I1=>b,
                O=>sig_159);
sigI_160 : and_2
      port map (I0=>a(160),
                I1=>b,
                O=>sig_160);
sigI_161 : and_2
      port map (I0=>a(161),
                I1=>b,
                O=>sig_161);				
sigI_162 : and_2
      port map (I0=>a(162),
                I1=>b,
                O=>sig_162);
xorI_162 : xor_2b
      port map (I0=>sig_162,
                I1=>c161_DUMMY,
                O=>xor_162);
xorI_161 : xor_2b
      port map (I0=>sig_161,
                I1=>c160_DUMMY,
                O=>xor_161);
xorI_160 : xor_2b
      port map (I0=>sig_160,
                I1=>c159_DUMMY,
                O=>xor_160);
xorI_159 : xor_2b
      port map (I0=>sig_159,
                I1=>c158_DUMMY,
                O=>xor_159);
xorI_158 : xor_2b
      port map (I0=>sig_158,
                I1=>c157_DUMMY,
                O=>xor_158);
xorI_157 : xor_2b
      port map (I0=>sig_157,
                I1=>c156_DUMMY,
                O=>xor_157);
xorI_156 : xor_2b
      port map (I0=>sig_156,
                I1=>c155_DUMMY,
                O=>xor_156);
xorI_155 : xor_2b
      port map (I0=>sig_155,
                I1=>c154_DUMMY,
                O=>xor_155);
xorI_154 : xor_2b
      port map (I0=>sig_154,
                I1=>c153_DUMMY,
                O=>xor_154);
xorI_153 : xor_2b
      port map (I0=>sig_153,
                I1=>c152_DUMMY,
                O=>xor_153);
xorI_152 : xor_2b
      port map (I0=>sig_152,
                I1=>c151_DUMMY,
                O=>xor_152);
xorI_151 : xor_2b
      port map (I0=>sig_151,
                I1=>c150_DUMMY,
                O=>xor_151);
xorI_150 : xor_2b
      port map (I0=>sig_150,
                I1=>c149_DUMMY,
                O=>xor_150);
xorI_149 : xor_2b
      port map (I0=>sig_149,
                I1=>c148_DUMMY,
                O=>xor_149);
xorI_148 : xor_2b
      port map (I0=>sig_148,
                I1=>c147_DUMMY,
                O=>xor_148);
xorI_147 : xor_2b
      port map (I0=>sig_147,
                I1=>c146_DUMMY,
                O=>xor_147);
xorI_146 : xor_2b
      port map (I0=>sig_146,
                I1=>c145_DUMMY,
                O=>xor_146);
xorI_145 : xor_2b
      port map (I0=>sig_145,
                I1=>c144_DUMMY,
                O=>xor_145);
xorI_144 : xor_2b
      port map (I0=>sig_144,
                I1=>c143_DUMMY,
                O=>xor_144);
xorI_143 : xor_2b
      port map (I0=>sig_143,
                I1=>c142_DUMMY,
                O=>xor_143);
xorI_142 : xor_2b
      port map (I0=>sig_142,
                I1=>c141_DUMMY,
                O=>xor_142);
xorI_141 : xor_2b
      port map (I0=>sig_141,
                I1=>c140_DUMMY,
                O=>xor_141);
xorI_140 : xor_2b
      port map (I0=>sig_140,
                I1=>c139_DUMMY,
                O=>xor_140);
xorI_139 : xor_2b
      port map (I0=>sig_139,
                I1=>c138_DUMMY,
                O=>xor_139);
xorI_138 : xor_2b
      port map (I0=>sig_138,
                I1=>c137_DUMMY,
                O=>xor_138);
xorI_137 : xor_2b
      port map (I0=>sig_137,
                I1=>c136_DUMMY,
                O=>xor_137);
xorI_136 : xor_2b
      port map (I0=>sig_136,
                I1=>c135_DUMMY,
                O=>xor_136);
xorI_135 : xor_2b
      port map (I0=>sig_135,
                I1=>c134_DUMMY,
                O=>xor_135);
xorI_134 : xor_2b
      port map (I0=>sig_134,
                I1=>c133_DUMMY,
                O=>xor_134);
xorI_133 : xor_2b
      port map (I0=>sig_133,
                I1=>c132_DUMMY,
                O=>xor_133);
xorI_132 : xor_2b
      port map (I0=>sig_132,
                I1=>c131_DUMMY,
                O=>xor_132);
xorI_131 : xor_2b
      port map (I0=>sig_131,
                I1=>c130_DUMMY,
                O=>xor_131);
xorI_130 : xor_2b
      port map (I0=>sig_130,
                I1=>c129_DUMMY,
                O=>xor_130);
xorI_129 : xor_2b
      port map (I0=>sig_129,
                I1=>c128_DUMMY,
                O=>xor_129);
xorI_128 : xor_2b
      port map (I0=>sig_128,
                I1=>c127_DUMMY,
                O=>xor_128);
xorI_127 : xor_2b
      port map (I0=>sig_127,
                I1=>c126_DUMMY,
                O=>xor_127);
xorI_126 : xor_2b
      port map (I0=>sig_126,
                I1=>c125_DUMMY,
                O=>xor_126);
xorI_125 : xor_2b
      port map (I0=>sig_125,
                I1=>c124_DUMMY,
                O=>xor_125);
xorI_124 : xor_2b
      port map (I0=>sig_124,
                I1=>c123_DUMMY,
                O=>xor_124);
xorI_123 : xor_2b
      port map (I0=>sig_123,
                I1=>c122_DUMMY,
                O=>xor_123);
xorI_122 : xor_2b
      port map (I0=>sig_122,
                I1=>c121_DUMMY,
                O=>xor_122);
xorI_121 : xor_2b
      port map (I0=>sig_121,
                I1=>c120_DUMMY,
                O=>xor_121);
xorI_120 : xor_2b
      port map (I0=>sig_120,
                I1=>c119_DUMMY,
                O=>xor_120);
xorI_119 : xor_2b
      port map (I0=>sig_119,
                I1=>c118_DUMMY,
                O=>xor_119);
xorI_118 : xor_2b
      port map (I0=>sig_118,
                I1=>c117_DUMMY,
                O=>xor_118);
xorI_117 : xor_2b
      port map (I0=>sig_117,
                I1=>c116_DUMMY,
                O=>xor_117);
xorI_116 : xor_2b
      port map (I0=>sig_116,
                I1=>c115_DUMMY,
                O=>xor_116);
xorI_115 : xor_2b
      port map (I0=>sig_115,
                I1=>c114_DUMMY,
                O=>xor_115);
xorI_114 : xor_2b
      port map (I0=>sig_114,
                I1=>c113_DUMMY,
                O=>xor_114);
xorI_113 : xor_2b
      port map (I0=>sig_113,
                I1=>c112_DUMMY,
                O=>xor_113);
xorI_112 : xor_2b
      port map (I0=>sig_112,
                I1=>c111_DUMMY,
                O=>xor_112);
xorI_111 : xor_2b
      port map (I0=>sig_111,
                I1=>c110_DUMMY,
                O=>xor_111);
xorI_110 : xor_2b
      port map (I0=>sig_110,
                I1=>c109_DUMMY,
                O=>xor_110);
xorI_109 : xor_2b
      port map (I0=>sig_109,
                I1=>c108_DUMMY,
                O=>xor_109);
xorI_108 : xor_2b
      port map (I0=>sig_108,
                I1=>c107_DUMMY,
                O=>xor_108);
xorI_107 : xor_2b
      port map (I0=>sig_107,
                I1=>c106_DUMMY,
                O=>xor_107);
xorI_106 : xor_2b
      port map (I0=>sig_106,
                I1=>c105_DUMMY,
                O=>xor_106);
xorI_105 : xor_2b
      port map (I0=>sig_105,
                I1=>c104_DUMMY,
                O=>xor_105);
xorI_104 : xor_2b
      port map (I0=>sig_104,
                I1=>c103_DUMMY,
                O=>xor_104);
xorI_103 : xor_2b
      port map (I0=>sig_103,
                I1=>c102_DUMMY,
                O=>xor_103);
xorI_102 : xor_2b
      port map (I0=>sig_102,
                I1=>c101_DUMMY,
                O=>xor_102);
xorI_101 : xor_2b
      port map (I0=>sig_101,
                I1=>c100_DUMMY,
                O=>xor_101);
xorI_100 : xor_2b
      port map (I0=>sig_100,
                I1=>c99_DUMMY,
                O=>xor_100);
xorI_99 : xor_2b
      port map (I0=>sig_99,
                I1=>c98_DUMMY,
                O=>xor_99);
xorI_98 : xor_2b
      port map (I0=>sig_98,
                I1=>c97_DUMMY,
                O=>xor_98);
xorI_97 : xor_2b
      port map (I0=>sig_97,
                I1=>c96_DUMMY,
                O=>xor_97);
xorI_96 : xor_2b
      port map (I0=>sig_96,
                I1=>c95_DUMMY,
                O=>xor_96);
xorI_95 : xor_2b
      port map (I0=>sig_95,
                I1=>c94_DUMMY,
                O=>xor_95);
xorI_94 : xor_2b
      port map (I0=>sig_94,
                I1=>c93_DUMMY,
                O=>xor_94);
xorI_93 : xor_2b
      port map (I0=>sig_93,
                I1=>c92_DUMMY,
                O=>xor_93);
xorI_92 : xor_2b
      port map (I0=>sig_92,
                I1=>c91_DUMMY,
                O=>xor_92);
xorI_91 : xor_2b
      port map (I0=>sig_91,
                I1=>c90_DUMMY,
                O=>xor_91);
xorI_90 : xor_2b
      port map (I0=>sig_90,
                I1=>c89_DUMMY,
                O=>xor_90);
xorI_89 : xor_2b
      port map (I0=>sig_89,
                I1=>c88_DUMMY,
                O=>xor_89);
xorI_88 : xor_2b
      port map (I0=>sig_88,
                I1=>c87_DUMMY,
                O=>xor_88);
xorI_87 : xor_2b
      port map (I0=>sig_87,
                I1=>c86_DUMMY,
                O=>xor_87);				
xorI_86 : xor_2b
      port map (I0=>sig_86,
                I1=>c85_DUMMY,
                O=>xor_86);
xorI_85 : xor_2b
      port map (I0=>sig_85,
                I1=>c84_DUMMY,
                O=>xor_85);	
xorI_84 : xor_2b
      port map (I0=>sig_84,
                I1=>c83_DUMMY,
                O=>xor_84);
xorI_83 : xor_2b
      port map (I0=>sig_83,
                I1=>c82_DUMMY,
                O=>xor_83);
xorI_82 : xor_2b
      port map (I0=>sig_82,
                I1=>c81_DUMMY,
                O=>xor_82);
xorI_81 : xor_2b
      port map (I0=>sig_81,
                I1=>c80_DUMMY,
                O=>xor_81);
xorI_80 : xor_2b
      port map (I0=>sig_80,
                I1=>c79_DUMMY,
                O=>xor_80);
xorI_79 : xor_2b
      port map (I0=>sig_79,
                I1=>c78_DUMMY,
                O=>xor_79);
xorI_78 : xor_2b
      port map (I0=>sig_78,
                I1=>c77_DUMMY,
                O=>xor_78);
xorI_77 : xor_2b
      port map (I0=>sig_77,
                I1=>c76_DUMMY,
                O=>xor_77);
xorI_76 : xor_2b
      port map (I0=>sig_76,
                I1=>c75_DUMMY,
                O=>xor_76);
xorI_75 : xor_2b
      port map (I0=>sig_75,
                I1=>c74_DUMMY,
                O=>xor_75);
xorI_74 : xor_2b
      port map (I0=>sig_74,
                I1=>c73_DUMMY,
                O=>xor_74);
xorI_73 : xor_2b
      port map (I0=>sig_73,
                I1=>c72_DUMMY,
                O=>xor_73);
xorI_72 : xor_2b
      port map (I0=>sig_72,
                I1=>c71_DUMMY,
                O=>xor_72);
xorI_71 : xor_2b
      port map (I0=>sig_71,
                I1=>c70_DUMMY,
                O=>xor_71);
xorI_70 : xor_2b
      port map (I0=>sig_70,
                I1=>c69_DUMMY,
                O=>xor_70);
xorI_69 : xor_2b
      port map (I0=>sig_69,
                I1=>c68_DUMMY,
                O=>xor_69);
xorI_68 : xor_2b
      port map (I0=>sig_68,
                I1=>c67_DUMMY,
                O=>xor_68);
xorI_67 : xor_2b
      port map (I0=>sig_67,
                I1=>c66_DUMMY,
                O=>xor_67);
xorI_66 : xor_2b
      port map (I0=>sig_66,
                I1=>c65_DUMMY,
                O=>xor_66);
xorI_65 : xor_2b
      port map (I0=>sig_65,
                I1=>c64_DUMMY,
                O=>xor_65);
xorI_64 : xor_2b
      port map (I0=>sig_64,
                I1=>c63_DUMMY,
                O=>xor_64);
xorI_63 : xor_2b
      port map (I0=>sig_63,
                I1=>c62_DUMMY,
                O=>xor_63);
xorI_62 : xor_2b
      port map (I0=>sig_62,
                I1=>c61_DUMMY,
                O=>xor_62);	
xorI_61 : xor_2b
      port map (I0=>sig_61,
                I1=>c60_DUMMY,
                O=>xor_61);
xorI_60 : xor_2b
      port map (I0=>sig_60,
                I1=>c59_DUMMY,
                O=>xor_60);
xorI_59 : xor_2b
      port map (I0=>sig_59,
                I1=>c58_DUMMY,
                O=>xor_59);
xorI_58 : xor_2b
      port map (I0=>sig_58,
                I1=>c57_DUMMY,
                O=>xor_58);
xorI_57 : xor_2b
      port map (I0=>sig_57,
                I1=>c56_DUMMY,
                O=>xor_57);
xorI_56 : xor_2b
      port map (I0=>sig_56,
                I1=>c55_DUMMY,
                O=>xor_56);
xorI_55 : xor_2b
      port map (I0=>sig_55,
                I1=>c54_DUMMY,
                O=>xor_55);
xorI_54 : xor_2b
      port map (I0=>sig_54,
                I1=>c53_DUMMY,
                O=>xor_54);
xorI_53 : xor_2b
      port map (I0=>sig_53,
                I1=>c52_DUMMY,
                O=>xor_53);
xorI_52 : xor_2b
      port map (I0=>sig_52,
                I1=>c51_DUMMY,
                O=>xor_52);
xorI_51 : xor_2b
      port map (I0=>sig_51,
                I1=>c50_DUMMY,
                O=>xor_51);	
xorI_50 : xor_2b
      port map (I0=>sig_50,
                I1=>c49_DUMMY,
                O=>xor_50);
xorI_49 : xor_2b
      port map (I0=>sig_49,
                I1=>c48_DUMMY,
                O=>xor_49);
xorI_48 : xor_2b
      port map (I0=>sig_48,
                I1=>c47_DUMMY,
                O=>xor_48);	
xorI_47 : xor_2b
      port map (I0=>sig_47,
                I1=>c46_DUMMY,
                O=>xor_47);	
xorI_46 : xor_2b
      port map (I0=>sig_46,
                I1=>c45_DUMMY,
                O=>xor_46);	
xorI_45 : xor_2b
      port map (I0=>sig_45,
                I1=>c44_DUMMY,
                O=>xor_45);	
xorI_44 : xor_2b
      port map (I0=>sig_44,
                I1=>c44_DUMMY,
                O=>xor_44);	
xorI_43 : xor_2b
      port map (I0=>sig_43,
                I1=>c42_DUMMY,
                O=>xor_43);	
xorI_42 : xor_2b
      port map (I0=>sig_42,
                I1=>c41_DUMMY,
                O=>xor_42);	
xorI_41 : xor_2b
      port map (I0=>sig_41,
                I1=>c40_DUMMY,
                O=>xor_41);
xorI_40 : xor_2b
      port map (I0=>sig_40,
                I1=>c39_DUMMY,
                O=>xor_40);
xorI_39 : xor_2b
      port map (I0=>sig_39,
                I1=>c38_DUMMY,
                O=>xor_39);	
xorI_38 : xor_2b
      port map (I0=>sig_38,
                I1=>c37_DUMMY,
                O=>xor_38);	
xorI_37 : xor_2b
      port map (I0=>sig_37,
                I1=>c36_DUMMY,
                O=>xor_37);
xorI_36 : xor_2b
      port map (I0=>sig_36,
                I1=>c35_DUMMY,
                O=>xor_36);	
xorI_35 : xor_2b
      port map (I0=>sig_35,
                I1=>c34_DUMMY,
                O=>xor_35);
xorI_34 : xor_2b
      port map (I0=>sig_34,
                I1=>c33_DUMMY,
                O=>xor_34);	
xorI_33 : xor_2b
      port map (I0=>sig_33,
                I1=>c32_DUMMY,
                O=>xor_33);
xorI_32 : xor_2b
      port map (I0=>sig_32,
                I1=>c31_DUMMY,
                O=>xor_32);	
xorI_31 : xor_2b
      port map (I0=>sig_31,
                I1=>c30_DUMMY,
                O=>xor_31);
xorI_30 : xor_2b
      port map (I0=>sig_30,
                I1=>c29_DUMMY,
                O=>xor_30);
xorI_29 : xor_2b
      port map (I0=>sig_29,
                I1=>c28_DUMMY,
                O=>xor_29);
xorI_28 : xor_2b
      port map (I0=>sig_28,
                I1=>c27_DUMMY,
                O=>xor_28);
xorI_27 : xor_2b
      port map (I0=>sig_27,
                I1=>c26_DUMMY,
                O=>xor_27);
xorI_26 : xor_2b
      port map (I0=>sig_26,
                I1=>c25_DUMMY,
                O=>xor_26);
xorI_25 : xor_2b
      port map (I0=>sig_25,
                I1=>c24_DUMMY,
                O=>xor_25);
xorI_24 : xor_2b
      port map (I0=>sig_24,
                I1=>c23_DUMMY,
                O=>xor_24);
xorI_23 : xor_2b
      port map (I0=>sig_23,
                I1=>c23_DUMMY,
                O=>xor_23);
xorI_22 : xor_2b
      port map (I0=>sig_22,
                I1=>c21_DUMMY,
                O=>xor_22);
xorI_21 : xor_2b
      port map (I0=>sig_21,
                I1=>c20_DUMMY,
                O=>xor_21);
xorI_20 : xor_2b
      port map (I0=>sig_20,
                I1=>c19_DUMMY,
                O=>xor_20);
xorI_19 : xor_2b
      port map (I0=>sig_19,
                I1=>c18_DUMMY,
                O=>xor_19);
xorI_18 : xor_2b
      port map (I0=>sig_18,
                I1=>c17_DUMMY,
                O=>xor_18);	
xorI_17 : xor_2b
      port map (I0=>sig_17,
                I1=>c16_DUMMY,
                O=>xor_17);
xorI_16 : xor_2b
      port map (I0=>sig_16,
                I1=>c15_DUMMY,
                O=>xor_16);
xorI_15 : xor_2b
      port map (I0=>sig_15,
                I1=>c14_DUMMY,
                O=>xor_15);	
xorI_14 : xor_2b
      port map (I0=>sig_14,
                I1=>c13_DUMMY,
                O=>xor_14);
xorI_13 : xor_2b
      port map (I0=>sig_13,
                I1=>c12_DUMMY,
                O=>xor_13);
xorI_12 : xor_2b
      port map (I0=>sig_12,
                I1=>c11_DUMMY,
                O=>xor_12);
xorI_11 : xor_2b
      port map (I0=>sig_11,
                I1=>c10_DUMMY,
                O=>xor_11);
xorI_10 : xor_2b
      port map (I0=>sig_10,
                I1=>c9_DUMMY,
                O=>xor_10);
xorI_9 : xor_2b
      port map (I0=>sig_9,
                I1=>c8_DUMMY,
                O=>xor_9);
xorI_8 : xor_2b
      port map (I0=>sig_8,
                I1=>c7_DUMMY,
                O=>xor_8);
xorI_c6c162 : xor_2b
      port map (I0=>c6_DUMMY,
                I1=>c162_DUMMY,
                O=>xor_c6c162);				
xorI_7 : xor_2b
      port map (I0=>sig_7,
                I1=>xor_c6c162,
                O=>xor_7);
xorI_c5c162 : xor_2b
      port map (I0=>c5_DUMMY,
                I1=>c162_DUMMY,
                O=>xor_c5c162);
xorI_6 : xor_2b
      port map (I0=>sig_6,
                I1=>xor_c5c162,
                O=>xor_6);
xorI_5 : xor_2b
      port map (I0=>sig_5,
                I1=>c4_DUMMY,
                O=>xor_5);
xorI_4 : xor_2b
      port map (I0=>sig_4,
                I1=>c3_DUMMY,
                O=>xor_4);
xorI_c2c162 : xor_2b
      port map (I0=>c2_DUMMY,
                I1=>c162_DUMMY,
                O=>xor_c2c162);
xorI_3 : xor_2b
      port map (I0=>sig_3,
                I1=>xor_c2c162,
                O=>xor_3);
xorI_2 : xor_2b
      port map (I0=>sig_2,
                I1=>c1_DUMMY,
                O=>xor_2);
xorI_1 : xor_2b
      port map (I0=>sig_1,
                I1=>c0_DUMMY,
                O=>xor_1);
   
xorI_0 : xor_2b
      port map (I0=>sig_0,
                I1=>c162_DUMMY,
                O=>xor_0);				
				
   reg_162 : reg_dff
      port map (D=>xor_162,
                clk=>clk,
				reset=>reset,
                Q=>c162_DUMMY);
   
   reg_161 : reg_dff
      port map (D=>xor_161,
                clk=>clk,
				reset=>reset,
                Q=>c161_DUMMY);
   
   reg_160 : reg_dff
      port map (D=>xor_160,
                clk=>clk,
				reset=>reset,
                Q=>c160_DUMMY);
   
   reg_159 : reg_dff
      port map (D=>xor_159,
	            clk=>clk,
                reset=>reset,
                Q=>c159_DUMMY);
   reg_158 : reg_dff
      port map (D=>xor_158,
                clk=>clk,
				reset=>reset,
                Q=>c158_DUMMY);
   
   reg_157 : reg_dff
      port map (D=>xor_157,
                clk=>clk,
				reset=>reset,
                Q=>c157_DUMMY);
   
   reg_156 : reg_dff
      port map (D=>xor_156,
                clk=>clk,
				reset=>reset,
                Q=>c156_DUMMY);
   
   reg_155 : reg_dff
      port map (D=>xor_155,
	            clk=>clk,
                reset=>reset,
                Q=>c155_DUMMY);
   
   reg_154 : reg_dff
      port map (D=>xor_154,
                clk=>clk,
				reset=>reset,
                Q=>c154_DUMMY);				
   
   reg_153 : reg_dff
      port map (D=>xor_153,
                clk=>clk,
				reset=>reset,
                Q=>c153_DUMMY);
   reg_152 : reg_dff
      port map (D=>xor_152,
                clk=>clk,
				reset=>reset,
                Q=>c152_DUMMY);
   
   reg_151 : reg_dff
      port map (D=>xor_151,
                clk=>clk,
				reset=>reset,
                Q=>c151_DUMMY);
   
   reg_150 : reg_dff
      port map (D=>xor_150,
                clk=>clk,
				reset=>reset,
                Q=>c150_DUMMY);
   
   reg_149 : reg_dff
      port map (D=>xor_149,
	            clk=>clk,
                reset=>reset,
                Q=>c149_DUMMY);
   
   reg_148 : reg_dff
      port map (D=>xor_148,
                clk=>clk,
				reset=>reset,
                Q=>c148_DUMMY);
   reg_147 : reg_dff
      port map (D=>xor_147,
                clk=>clk,
				reset=>reset,
                Q=>c147_DUMMY);
   
   reg_146 : reg_dff
      port map (D=>xor_146,
                clk=>clk,
				reset=>reset,
                Q=>c146_DUMMY);
   
   reg_145 : reg_dff
      port map (D=>xor_145,
                clk=>clk,
				reset=>reset,
                Q=>c145_DUMMY);
   
   reg_144 : reg_dff
      port map (D=>xor_144,
	            clk=>clk,
                reset=>reset,
                Q=>c144_DUMMY);
   
   reg_143 : reg_dff
      port map (D=>xor_143,
                clk=>clk,
				reset=>reset,
                Q=>c143_DUMMY);
   reg_142 : reg_dff
      port map (D=>xor_142,
                clk=>clk,
				reset=>reset,
                Q=>c142_DUMMY);
   
   reg_141 : reg_dff
      port map (D=>xor_141,
                clk=>clk,
				reset=>reset,
                Q=>c141_DUMMY);
   
   reg_140 : reg_dff
      port map (D=>xor_140,
                clk=>clk,
				reset=>reset,
                Q=>c140_DUMMY);
   
   reg_139 : reg_dff
      port map (D=>xor_139,
	            clk=>clk,
                reset=>reset,
                Q=>c139_DUMMY);
   
   reg_138 : reg_dff
      port map (D=>xor_138,
                clk=>clk,
				reset=>reset,
                Q=>c138_DUMMY);
   reg_137 : reg_dff
      port map (D=>xor_137,
                clk=>clk,
				reset=>reset,
                Q=>c137_DUMMY);
   
   reg_136 : reg_dff
      port map (D=>xor_136,
                clk=>clk,
				reset=>reset,
                Q=>c136_DUMMY);
   
   reg_135 : reg_dff
      port map (D=>xor_135,
                clk=>clk,
				reset=>reset,
                Q=>c135_DUMMY);
   
   reg_134 : reg_dff
      port map (D=>xor_134,
	            clk=>clk,
                reset=>reset,
                Q=>c134_DUMMY);
   
   reg_133 : reg_dff
      port map (D=>xor_133,
                clk=>clk,
				reset=>reset,
                Q=>c133_DUMMY);
   reg_132 : reg_dff
      port map (D=>xor_132,
                clk=>clk,
				reset=>reset,
                Q=>c132_DUMMY);
   
   reg_131 : reg_dff
      port map (D=>xor_131,
                clk=>clk,
				reset=>reset,
                Q=>c131_DUMMY);
   
   reg_130 : reg_dff
      port map (D=>xor_130,
                clk=>clk,
				reset=>reset,
                Q=>c130_DUMMY);
   
   reg_129 : reg_dff
      port map (D=>xor_129,
	            clk=>clk,
                reset=>reset,
                Q=>c129_DUMMY);
   
   reg_128 : reg_dff
      port map (D=>xor_128,
                clk=>clk,
				reset=>reset,
                Q=>c128_DUMMY);	
   reg_127 : reg_dff
      port map (D=>xor_127,
                clk=>clk,
				reset=>reset,
                Q=>c127_DUMMY);
   
   reg_126 : reg_dff
      port map (D=>xor_126,
                clk=>clk,
				reset=>reset,
                Q=>c126_DUMMY);
   
   reg_125 : reg_dff
      port map (D=>xor_125,
                clk=>clk,
				reset=>reset,
                Q=>c125_DUMMY);
   
   reg_124 : reg_dff
      port map (D=>xor_124,
	            clk=>clk,
                reset=>reset,
                Q=>c124_DUMMY);
   
   reg_123 : reg_dff
      port map (D=>xor_123,
                clk=>clk,
				reset=>reset,
                Q=>c123_DUMMY);	
   reg_122 : reg_dff
      port map (D=>xor_122,
                clk=>clk,
				reset=>reset,
                Q=>c122_DUMMY);
   
   reg_121 : reg_dff
      port map (D=>xor_121,
                clk=>clk,
				reset=>reset,
                Q=>c121_DUMMY);
   
   reg_120 : reg_dff
      port map (D=>xor_120,
                clk=>clk,
				reset=>reset,
                Q=>c120_DUMMY);
   
   reg_119 : reg_dff
      port map (D=>xor_119,
	            clk=>clk,
                reset=>reset,
                Q=>c119_DUMMY);
   
   reg_118 : reg_dff
      port map (D=>xor_118,
                clk=>clk,
				reset=>reset,
                Q=>c118_DUMMY);	
   reg_117 : reg_dff
      port map (D=>xor_117,
                clk=>clk,
				reset=>reset,
                Q=>c117_DUMMY);
   
   reg_116 : reg_dff
      port map (D=>xor_116,
                clk=>clk,
				reset=>reset,
                Q=>c116_DUMMY);
   
   reg_115 : reg_dff
      port map (D=>xor_115,
                clk=>clk,
				reset=>reset,
                Q=>c115_DUMMY);
   
   reg_114 : reg_dff
      port map (D=>xor_114,
	            clk=>clk,
                reset=>reset,
                Q=>c114_DUMMY);
   
   reg_113 : reg_dff
      port map (D=>xor_113,
                clk=>clk,
				reset=>reset,
                Q=>c113_DUMMY);
   reg_112 : reg_dff
      port map (D=>xor_112,
                clk=>clk,
				reset=>reset,
                Q=>c112_DUMMY);
   
   reg_111 : reg_dff
      port map (D=>xor_111,
                clk=>clk,
				reset=>reset,
                Q=>c111_DUMMY);
   
   reg_110 : reg_dff
      port map (D=>xor_110,
                clk=>clk,
				reset=>reset,
                Q=>c110_DUMMY);
   
   reg_109 : reg_dff
      port map (D=>xor_109,
	            clk=>clk,
                reset=>reset,
                Q=>c109_DUMMY);
   
   reg_108 : reg_dff
      port map (D=>xor_108,
                clk=>clk,
				reset=>reset,
                Q=>c108_DUMMY);
   reg_107 : reg_dff
      port map (D=>xor_107,
                clk=>clk,
				reset=>reset,
                Q=>c107_DUMMY);
   
   reg_106 : reg_dff
      port map (D=>xor_106,
                clk=>clk,
				reset=>reset,
                Q=>c106_DUMMY);
   
   reg_105 : reg_dff
      port map (D=>xor_105,
                clk=>clk,
				reset=>reset,
                Q=>c105_DUMMY);
   
   reg_104 : reg_dff
      port map (D=>xor_104,
	            clk=>clk,
                reset=>reset,
                Q=>c104_DUMMY);
   
   reg_103 : reg_dff
      port map (D=>xor_103,
                clk=>clk,
				reset=>reset,
                Q=>c103_DUMMY);
   reg_102 : reg_dff
      port map (D=>xor_102,
                clk=>clk,
				reset=>reset,
                Q=>c102_DUMMY);
   
   reg_101 : reg_dff
      port map (D=>xor_101,
                clk=>clk,
				reset=>reset,
                Q=>c101_DUMMY);
   
   reg_100 : reg_dff
      port map (D=>xor_100,
                clk=>clk,
				reset=>reset,
                Q=>c100_DUMMY);
   
   reg_99 : reg_dff
      port map (D=>xor_99,
	            clk=>clk,
                reset=>reset,
                Q=>c99_DUMMY);
   
   reg_98 : reg_dff
      port map (D=>xor_98,
                clk=>clk,
				reset=>reset,
                Q=>c98_DUMMY);
   reg_97 : reg_dff
      port map (D=>xor_97,
                clk=>clk,
				reset=>reset,
                Q=>c97_DUMMY);
   
   reg_96 : reg_dff
      port map (D=>xor_96,
                clk=>clk,
				reset=>reset,
                Q=>c96_DUMMY);
   
   reg_95 : reg_dff
      port map (D=>xor_95,
                clk=>clk,
				reset=>reset,
                Q=>c95_DUMMY);
   
   reg_94 : reg_dff
      port map (D=>xor_94,
	            clk=>clk,
                reset=>reset,
                Q=>c94_DUMMY);
   
   reg_93 : reg_dff
      port map (D=>xor_93,
                clk=>clk,
				reset=>reset,
                Q=>c93_DUMMY);
   reg_92 : reg_dff
      port map (D=>xor_92,
                clk=>clk,
				reset=>reset,
                Q=>c92_DUMMY);
   
   reg_91 : reg_dff
      port map (D=>xor_91,
                clk=>clk,
				reset=>reset,
                Q=>c91_DUMMY);
   
   reg_90 : reg_dff
      port map (D=>xor_90,
                clk=>clk,
				reset=>reset,
                Q=>c90_DUMMY);
   
   reg_89 : reg_dff
      port map (D=>xor_89,
	            clk=>clk,
                reset=>reset,
                Q=>c89_DUMMY);
   
   reg_88 : reg_dff
      port map (D=>xor_88,
                clk=>clk,
				reset=>reset,
                Q=>c88_DUMMY);
   reg_87 : reg_dff
      port map (D=>xor_87,
                clk=>clk,
				reset=>reset,
                Q=>c87_DUMMY);
   
   reg_86 : reg_dff
      port map (D=>xor_86,
                clk=>clk,
				reset=>reset,
                Q=>c86_DUMMY);
   
   reg_85 : reg_dff
      port map (D=>xor_85,
                clk=>clk,
				reset=>reset,
                Q=>c85_DUMMY);
   
   reg_84 : reg_dff
      port map (D=>xor_84,
	            clk=>clk,
                reset=>reset,
                Q=>c84_DUMMY);
   
   reg_83 : reg_dff
      port map (D=>xor_83,
                clk=>clk,
				reset=>reset,
                Q=>c83_DUMMY);
   reg_82 : reg_dff
      port map (D=>xor_82,
                clk=>clk,
				reset=>reset,
                Q=>c82_DUMMY);
   
   reg_81 : reg_dff
      port map (D=>xor_81,
                clk=>clk,
				reset=>reset,
                Q=>c81_DUMMY);
   
   reg_80 : reg_dff
      port map (D=>xor_80,
                clk=>clk,
				reset=>reset,
                Q=>c80_DUMMY);
   
   reg_79 : reg_dff
      port map (D=>xor_79,
	            clk=>clk,
                reset=>reset,
                Q=>c79_DUMMY);
   
   reg_78 : reg_dff
      port map (D=>xor_78,
                clk=>clk,
				reset=>reset,
                Q=>c78_DUMMY);
   reg_77 : reg_dff
      port map (D=>xor_77,
                clk=>clk,
				reset=>reset,
                Q=>c77_DUMMY);
   
   reg_76 : reg_dff
      port map (D=>xor_76,
                clk=>clk,
				reset=>reset,
                Q=>c76_DUMMY);
   
   reg_75 : reg_dff
      port map (D=>xor_75,
                clk=>clk,
				reset=>reset,
                Q=>c75_DUMMY);
   
   reg_74 : reg_dff
      port map (D=>xor_74,
	            clk=>clk,
                reset=>reset,
                Q=>c74_DUMMY);
   
   reg_73 : reg_dff
      port map (D=>xor_73,
                clk=>clk,
				reset=>reset,
                Q=>c73_DUMMY);
   reg_72 : reg_dff
      port map (D=>xor_72,
                clk=>clk,
				reset=>reset,
                Q=>c72_DUMMY);
   
   reg_71 : reg_dff
      port map (D=>xor_71,
                clk=>clk,
				reset=>reset,
                Q=>c71_DUMMY);
   
   reg_70 : reg_dff
      port map (D=>xor_70,
                clk=>clk,
				reset=>reset,
                Q=>c70_DUMMY);
   
   reg_69 : reg_dff
      port map (D=>xor_69,
	            clk=>clk,
                reset=>reset,
                Q=>c69_DUMMY);
   
   reg_68 : reg_dff
      port map (D=>xor_68,
                clk=>clk,
				reset=>reset,
                Q=>c68_DUMMY);
   reg_67 : reg_dff
      port map (D=>xor_67,
                clk=>clk,
				reset=>reset,
                Q=>c67_DUMMY);
   
   reg_66 : reg_dff
      port map (D=>xor_66,
                clk=>clk,
				reset=>reset,
                Q=>c66_DUMMY);
   
   reg_65 : reg_dff
      port map (D=>xor_65,
                clk=>clk,
				reset=>reset,
                Q=>c65_DUMMY);
   
   reg_64 : reg_dff
      port map (D=>xor_64,
	            clk=>clk,
                reset=>reset,
                Q=>c64_DUMMY);
   
   reg_63 : reg_dff
      port map (D=>xor_63,
                clk=>clk,
				reset=>reset,
                Q=>c63_DUMMY);
   reg_62 : reg_dff
      port map (D=>xor_62,
                clk=>clk,
				reset=>reset,
                Q=>c62_DUMMY);
   
   reg_61 : reg_dff
      port map (D=>xor_61,
                clk=>clk,
				reset=>reset,
                Q=>c61_DUMMY);
   
   reg_60 : reg_dff
      port map (D=>xor_60,
                clk=>clk,
				reset=>reset,
                Q=>c60_DUMMY);
   
   reg_59 : reg_dff
      port map (D=>xor_59,
	            clk=>clk,
                reset=>reset,
                Q=>c59_DUMMY);
   
   reg_58 : reg_dff
      port map (D=>xor_58,
                clk=>clk,
				reset=>reset,
                Q=>c58_DUMMY);
   reg_57 : reg_dff
      port map (D=>xor_57,
                clk=>clk,
				reset=>reset,
                Q=>c57_DUMMY);
   
   reg_56 : reg_dff
      port map (D=>xor_56,
                clk=>clk,
				reset=>reset,
                Q=>c56_DUMMY);
   
   reg_55 : reg_dff
      port map (D=>xor_55,
                clk=>clk,
				reset=>reset,
                Q=>c55_DUMMY);
   
   reg_54 : reg_dff
      port map (D=>xor_54,
	            clk=>clk,
                reset=>reset,
                Q=>c54_DUMMY);
   
   reg_53 : reg_dff
      port map (D=>xor_53,
                clk=>clk,
				reset=>reset,
                Q=>c53_DUMMY);
 
   reg_52 : reg_dff
      port map (D=>xor_52,
                clk=>clk,
				reset=>reset,
                Q=>c52_DUMMY);
   
   reg_51 : reg_dff
      port map (D=>xor_51,
                clk=>clk,
				reset=>reset,
                Q=>c51_DUMMY);
   
   reg_50 : reg_dff
      port map (D=>xor_50,
	            clk=>clk,
                reset=>reset,
                Q=>c50_DUMMY);
   
   reg_49 : reg_dff
      port map (D=>xor_49,
                clk=>clk,
				reset=>reset,
                Q=>c49_DUMMY);
 
   reg_48 : reg_dff
      port map (D=>xor_48,
                clk=>clk,
				reset=>reset,
                Q=>c48_DUMMY);
   
   reg_47 : reg_dff
      port map (D=>xor_47,
                clk=>clk,
				reset=>reset,
                Q=>c47_DUMMY);
   
   reg_46 : reg_dff
      port map (D=>xor_46,
	            clk=>clk,
                reset=>reset,
                Q=>c46_DUMMY);
   
   reg_45 : reg_dff
      port map (D=>xor_45,
                clk=>clk,
				reset=>reset,
                Q=>c45_DUMMY);
 
   reg_44 : reg_dff
      port map (D=>xor_44,
                clk=>clk,
				reset=>reset,
                Q=>c44_DUMMY);
   
   reg_43 : reg_dff
      port map (D=>xor_43,
                clk=>clk,
				reset=>reset,
                Q=>c43_DUMMY);
   
   reg_42 : reg_dff
      port map (D=>xor_42,
	            clk=>clk,
                reset=>reset,
                Q=>c42_DUMMY);
   
   reg_41 : reg_dff
      port map (D=>xor_41,
                clk=>clk,
				reset=>reset,
                Q=>c41_DUMMY);
 
   reg_40 : reg_dff
      port map (D=>xor_40,
                clk=>clk,
				reset=>reset,
                Q=>c40_DUMMY);
   
   reg_39 : reg_dff
      port map (D=>xor_39,
                clk=>clk,
				reset=>reset,
                Q=>c39_DUMMY);
   
   reg_38 : reg_dff
      port map (D=>xor_38,
	            clk=>clk,
                reset=>reset,
                Q=>c38_DUMMY);
   
   reg_37 : reg_dff
      port map (D=>xor_37,
                clk=>clk,
				reset=>reset,
                Q=>c37_DUMMY);
 
   reg_36 : reg_dff
      port map (D=>xor_36,
                clk=>clk,
				reset=>reset,
                Q=>c36_DUMMY);
   
   reg_35 : reg_dff
      port map (D=>xor_35,
                clk=>clk,
				reset=>reset,
                Q=>c35_DUMMY);
   
   reg_34 : reg_dff
      port map (D=>xor_34,
	            clk=>clk,
                reset=>reset,
                Q=>c34_DUMMY);
   
   reg_33 : reg_dff
      port map (D=>xor_33,
                clk=>clk,
				reset=>reset,
                Q=>c33_DUMMY);
 
   reg_32 : reg_dff
      port map (D=>xor_32,
                clk=>clk,
				reset=>reset,
                Q=>c32_DUMMY);
   
   reg_31 : reg_dff
      port map (D=>xor_31,
                clk=>clk,
				reset=>reset,
                Q=>c31_DUMMY);
   
   reg_30 : reg_dff
      port map (D=>xor_30,
	            clk=>clk,
                reset=>reset,
                Q=>c30_DUMMY);
   
   reg_29 : reg_dff
      port map (D=>xor_29,
                clk=>clk,
				reset=>reset,
                Q=>c29_DUMMY);
 
   reg_28 : reg_dff
      port map (D=>xor_28,
                clk=>clk,
				reset=>reset,
                Q=>c28_DUMMY);
   
   reg_27 : reg_dff
      port map (D=>xor_27,
                clk=>clk,
				reset=>reset,
                Q=>c27_DUMMY);
   
   reg_26 : reg_dff
      port map (D=>xor_26,
	            clk=>clk,
                reset=>reset,
                Q=>c26_DUMMY);
   
   reg_25 : reg_dff
      port map (D=>xor_25,
                clk=>clk,
				reset=>reset,
                Q=>c25_DUMMY);
 
   reg_24 : reg_dff
      port map (D=>xor_24,
                clk=>clk,
				reset=>reset,
                Q=>c24_DUMMY);
   
   reg_23 : reg_dff
      port map (D=>xor_23,
                clk=>clk,
				reset=>reset,
                Q=>c23_DUMMY);
   
   reg_22 : reg_dff
      port map (D=>xor_22,
	            clk=>clk,
                reset=>reset,
                Q=>c22_DUMMY);
   
   reg_21 : reg_dff
      port map (D=>xor_21,
                clk=>clk,
				reset=>reset,
                Q=>c21_DUMMY);
 
   reg_20 : reg_dff
      port map (D=>xor_20,
                clk=>clk,
				reset=>reset,
                Q=>c20_DUMMY);
   
   reg_19 : reg_dff
      port map (D=>xor_19,
                clk=>clk,
				reset=>reset,
                Q=>c19_DUMMY);
   
   reg_18 : reg_dff
      port map (D=>xor_18,
	            clk=>clk,
                reset=>reset,
                Q=>c18_DUMMY);
   
   reg_17 : reg_dff
      port map (D=>xor_17,
                clk=>clk,
				reset=>reset,
                Q=>c17_DUMMY);
 
   reg_16 : reg_dff
      port map (D=>xor_16,
                clk=>clk,
				reset=>reset,
                Q=>c16_DUMMY);
   
   reg_15 : reg_dff
      port map (D=>xor_15,
                clk=>clk,
				reset=>reset,
                Q=>c15_DUMMY);
   
   reg_14 : reg_dff
      port map (D=>xor_14,
	            clk=>clk,
                reset=>reset,
                Q=>c14_DUMMY);
   
   reg_13 : reg_dff
      port map (D=>xor_13,
                clk=>clk,
				reset=>reset,
                Q=>c13_DUMMY);
 
   reg_12 : reg_dff
      port map (D=>xor_12,
                clk=>clk,
				reset=>reset,
                Q=>c12_DUMMY);
   
   reg_11 : reg_dff
      port map (D=>xor_11,
                clk=>clk,
				reset=>reset,
                Q=>c11_DUMMY);
   
   reg_10 : reg_dff
      port map (D=>xor_10,
	            clk=>clk,
                reset=>reset,
                Q=>c10_DUMMY);
   
   reg_9 : reg_dff
      port map (D=>xor_9,
                clk=>clk,
				reset=>reset,
                Q=>c9_DUMMY);
 
   reg_8 : reg_dff
      port map (D=>xor_8,
                clk=>clk,
				reset=>reset,
                Q=>c8_DUMMY);
   
   reg_7 : reg_dff
      port map (D=>xor_7,
                clk=>clk,
				reset=>reset,
                Q=>c7_DUMMY);
   
   reg_6 : reg_dff
      port map (D=>xor_6,
	            clk=>clk,
                reset=>reset,
                Q=>c6_DUMMY);
   
   reg_5 : reg_dff
      port map (D=>xor_5,
                clk=>clk,
				reset=>reset,
                Q=>c5_DUMMY);
  
   reg_4 : reg_dff
      port map (D=>xor_4,
                clk=>clk,
				reset=>reset,
                Q=>c4_DUMMY);
   
   reg_3 : reg_dff
      port map (D=>xor_3,
                clk=>clk,
				reset=>reset,
                Q=>c3_DUMMY);
   
   reg_2 : reg_dff
      port map (D=>xor_2,
                clk=>clk,
				reset=>reset,
                Q=>c2_DUMMY);
   
   reg_1 : reg_dff
      port map (D=>xor_1,
	            clk=>clk,
                reset=>reset,
                Q=>c1_DUMMY);
   
   reg_0 : reg_dff
      port map (D=>xor_0,
                clk=>clk,
				reset=>reset,
                Q=>c0_DUMMY);								
				
c(0) <= c0_DUMMY;				
c(1) <= c1_DUMMY;
c(2) <= c2_DUMMY;
c(3) <= c3_DUMMY;
c(4) <= c4_DUMMY;
c(5) <= c5_DUMMY;				
c(6) <= c6_DUMMY;
c(7) <= c7_DUMMY;
c(8) <= c8_DUMMY;
c(9) <= c9_DUMMY;
c(10) <= c10_DUMMY;				
c(11) <= c11_DUMMY;
c(12) <= c12_DUMMY;
c(13) <= c13_DUMMY;
c(14) <= c14_DUMMY;
c(15) <= c15_DUMMY;				
c(16) <= c16_DUMMY;
c(17) <= c17_DUMMY;
c(18) <= c18_DUMMY;
c(19) <= c19_DUMMY;
c(20) <= c20_DUMMY;				
c(21) <= c21_DUMMY;
c(22) <= c22_DUMMY;
c(23) <= c23_DUMMY;
c(24) <= c24_DUMMY;
c(25) <= c25_DUMMY;				
c(26) <= c26_DUMMY;
c(27) <= c27_DUMMY;
c(28) <= c28_DUMMY;
c(29) <= c29_DUMMY;
c(30) <= c30_DUMMY;				
c(31) <= c31_DUMMY;
c(32) <= c32_DUMMY;
c(33) <= c33_DUMMY;
c(34) <= c34_DUMMY;
c(35) <= c35_DUMMY;				
c(36) <= c36_DUMMY;
c(37) <= c37_DUMMY;
c(38) <= c38_DUMMY;
c(39) <= c39_DUMMY;
c(40) <= c40_DUMMY;				
c(41) <= c41_DUMMY;
c(42) <= c42_DUMMY;
c(43) <= c43_DUMMY;
c(44) <= c44_DUMMY;
c(45) <= c45_DUMMY;				
c(46) <= c46_DUMMY;
c(47) <= c47_DUMMY;
c(48) <= c48_DUMMY;
c(49) <= c49_DUMMY;
c(50) <= c50_DUMMY;				
c(51) <= c51_DUMMY;
c(52) <= c52_DUMMY;
c(53) <= c53_DUMMY;
c(54) <= c54_DUMMY;
c(55) <= c55_DUMMY;				
c(56) <= c56_DUMMY;
c(57) <= c57_DUMMY;
c(58) <= c58_DUMMY;
c(59) <= c59_DUMMY;
c(60) <= c60_DUMMY;				
c(61) <= c61_DUMMY;
c(62) <= c62_DUMMY;
c(63) <= c63_DUMMY;
c(64) <= c64_DUMMY;
c(65) <= c65_DUMMY;				
c(66) <= c66_DUMMY;
c(67) <= c67_DUMMY;
c(68) <= c68_DUMMY;
c(69) <= c69_DUMMY;
c(70) <= c70_DUMMY;				
c(71) <= c71_DUMMY;
c(72) <= c72_DUMMY;
c(73) <= c73_DUMMY;
c(74) <= c74_DUMMY;
c(75) <= c75_DUMMY;				
c(76) <= c76_DUMMY;
c(77) <= c77_DUMMY;
c(78) <= c78_DUMMY;
c(79) <= c79_DUMMY;
c(80) <= c80_DUMMY;				
c(81) <= c81_DUMMY;
c(82) <= c82_DUMMY;
c(83) <= c83_DUMMY;
c(84) <= c84_DUMMY;
c(85) <= c85_DUMMY;				
c(86) <= c86_DUMMY;
c(87) <= c87_DUMMY;
c(88) <= c88_DUMMY;
c(89) <= c89_DUMMY;
c(90) <= c90_DUMMY;				
c(91) <= c91_DUMMY;
c(92) <= c92_DUMMY;
c(93) <= c93_DUMMY;
c(94) <= c94_DUMMY;
c(95) <= c95_DUMMY;				
c(96) <= c96_DUMMY;
c(97) <= c97_DUMMY;
c(98) <= c98_DUMMY;
c(99) <= c99_DUMMY;
c(100) <= c100_DUMMY;				
c(101) <= c101_DUMMY;
c(102) <= c102_DUMMY;
c(103) <= c103_DUMMY;
c(104) <= c104_DUMMY;
c(105) <= c105_DUMMY;				
c(106) <= c106_DUMMY;
c(107) <= c107_DUMMY;
c(108) <= c108_DUMMY;
c(109) <= c109_DUMMY;
c(110) <= c110_DUMMY;				
c(111) <= c111_DUMMY;
c(112) <= c112_DUMMY;
c(113) <= c113_DUMMY;
c(114) <= c114_DUMMY;
c(115) <= c115_DUMMY;				
c(116) <= c116_DUMMY;
c(117) <= c117_DUMMY;
c(118) <= c118_DUMMY;
c(119) <= c119_DUMMY;
c(120) <= c120_DUMMY;				
c(121) <= c121_DUMMY;
c(122) <= c122_DUMMY;
c(123) <= c123_DUMMY;
c(124) <= c124_DUMMY;
c(125) <= c125_DUMMY;				
c(126) <= c126_DUMMY;
c(127) <= c127_DUMMY;
c(128) <= c128_DUMMY;
c(129) <= c129_DUMMY;
c(130) <= c130_DUMMY;				
c(131) <= c131_DUMMY;
c(132) <= c132_DUMMY;
c(133) <= c133_DUMMY;
c(134) <= c134_DUMMY;
c(135) <= c135_DUMMY;				
c(136) <= c136_DUMMY;
c(137) <= c137_DUMMY;
c(138) <= c138_DUMMY;
c(139) <= c139_DUMMY;
c(140) <= c140_DUMMY;				
c(141) <= c141_DUMMY;
c(142) <= c142_DUMMY;
c(143) <= c143_DUMMY;
c(144) <= c144_DUMMY;
c(145) <= c145_DUMMY;				
c(146) <= c146_DUMMY;
c(147) <= c147_DUMMY;
c(148) <= c148_DUMMY;
c(149) <= c149_DUMMY;
c(150) <= c150_DUMMY;				
c(151) <= c151_DUMMY;
c(152) <= c152_DUMMY;
c(153) <= c153_DUMMY;
c(154) <= c154_DUMMY;
c(155) <= c155_DUMMY;				
c(156) <= c156_DUMMY;
c(157) <= c157_DUMMY;
c(158) <= c158_DUMMY;
c(159) <= c159_DUMMY;
c(160) <= c160_DUMMY;
c(161) <= c161_DUMMY;
c(162) <= c162_DUMMY;					


end Behavioral;

